module top_module(input in,output out);
  not n(out,in);
endmodule
