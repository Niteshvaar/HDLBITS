module top_module ( input a, input b, output out );
    mod_a x(a,b,out);
endmodule
